library ieee;
library vunit_lib;
context vunit_lib.vunit_context; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity tb_counter is
  generic (runner_cfg : string);
end tb_counter;

architecture arch_tb_counter of tb_counter is
  component counter is
    port (
      key0: in std_logic;
      key3: in std_logic;
      counter_out: out std_logic_vector(3 downto 0)
    );
  end component;
  signal key0, key3: std_logic;
  signal counter_out: std_logic_vector(3 downto 0);

begin
  uut: counter port map(
    key0 => key0,
    key3 => key3,
    counter_out => counter_out
  );

  main: process
  procedure press_key0(constant x : std_logic) is
    begin
      key0 <= '0';
      wait for 50 ns; 
      key0 <= '1';
      wait for 45 ns; 
    end procedure;
  begin
    test_runner_setup(runner, runner_cfg);
    for j in 0 to 8 loop
      press_key0(key0);
      check_match(counter_out, (std_logic_vector(to_unsigned(j + 1, 4))));
    end loop;
    press_key0(key0);
    check_match(counter_out, "0000");
    test_runner_cleanup(runner); -- Simulation ends here
  end process;

end arch_tb_counter  ; -- arch_tb_counter 